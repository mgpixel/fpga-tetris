package types;

typedef enum logic [2:0] {
  EMPTY,
  CYAN,
  BLUE,
  ORANGE,
  YELLOW,
  GREEN,
  RED,
  MAGENTA
} block_color;

typedef enum logic [2:0] {
  I_CYAN,
  J_BLUE,
  L_ORANGE,
  O_YELLOW,
  P_GREEN,
  T_MAGENTA,
  Z_RED
} block_t;

typedef enum logic [1:0] {
  LEFT,
  RIGHT,
  DOWN
} direction;

typedef enum logic [1:0] {
  ROT_LEFT1,
  ROT_RIGHT1,
  ROT2,
  NORMAL
} orientation;

endpackage