// A pseudo random module to create blocks for the game. Most games have a bag of 7
// to be choosing from, this one just generates 1 block at a time. Holds the block index
// until a new one is needed.
module tetromino_generator
(
  input Clk,
  input Reset,
  input new_block,
  input logic [2:0] new_move,
  output logic [2:0] block_idx
);

logic [9:0] start = 10'd385;
logic [9:0] generated_bits = 10'd220;
logic [2:0] fair_idx;
logic [2:0] old_idx;

counter fair_counter(
  .Clk(Clk),
  .Reset(Reset || fair_idx > 3'd6),
  .load(new_block),
  .cur_val(fair_idx)
);

always_ff @(posedge Clk)
begin
  if (Reset) begin
    generated_bits <= generated_bits + start;
  end
  if (new_block)
    old_idx <= block_idx;
  generated_bits <= generated_bits + new_move + block_idx;
end

always_comb
begin
  block_idx = 3'd0;
  if (Reset)
    block_idx = generated_bits[5:3];
  else if (new_block) begin
    block_idx = generated_bits[2:0];
    if (block_idx > 3'd6 || block_idx == old_idx)
      block_idx = fair_idx;
  end
end

endmodule